module fpALU (

);
    
endmodule